module module_1;
endmodule

module module_2 #();
endmodule

module /* test */ module_3 #()(
    input clk_i
);
endmodule

module module_4 #()()(
    clk_i
);

input clk_i;
    module_1 i_module_1();
endmodule : module_4