package blub_pkg;

endpackage
