`include "include.svh"

module test;

logic d, q, clk_i, rst_ni;

`FF(q, d, '0)

endmodule